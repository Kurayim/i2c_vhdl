-- i2c
